* SPICE3 file created from sky130_fd_sc_hd__dfxtp_1.ext - technology: sky130A

.option scale=0.005u

.subckt sky130_fd_sc_hd__dfxtp_1 CLK D VGND VNB VPB VPWR Q
X0 a_975_413# a_193_47# a_891_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X1 VGND a_891_413# a_1059_315# VNB sky130_fd_pr__nfet_01v8 w=130 l=30
X2 a_561_413# a_27_47# a_466_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X3 a_891_413# a_27_47# a_634_159# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X4 a_466_413# a_193_47# a_381_47# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X5 a_381_47# D VPWR VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X6 a_634_159# a_466_413# VPWR VPB sky130_fd_pr__pfet_01v8 w=150 l=30
X7 a_634_159# a_466_413# VGND VNB sky130_fd_pr__nfet_01v8 w=128 l=30
X8 VGND a_1059_315# a_1017_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X9 VPWR a_891_413# a_1059_315# VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X10 VPWR a_634_159# a_561_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X11 Q a_1059_315# VPWR VPB sky130_fd_pr__pfet_01v8 w=200 l=30
X12 a_1017_47# a_27_47# a_891_413# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X13 a_891_413# a_193_47# a_634_159# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X14 VGND a_634_159# a_592_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X15 a_592_47# a_193_47# a_466_413# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X16 a_193_47# a_27_47# VGND VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X17 a_466_413# a_27_47# a_381_47# VNB sky130_fd_pr__nfet_01v8 w=72 l=30
X18 VGND CLK a_27_47# VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X19 VPWR CLK a_27_47# VPB sky130_fd_pr__pfet_01v8 w=128 l=30
X20 a_193_47# a_27_47# VPWR VPB sky130_fd_pr__pfet_01v8 w=128 l=30
X21 a_381_47# D VGND VNB sky130_fd_pr__nfet_01v8 w=84 l=30
X22 VPWR a_1059_315# a_975_413# VPB sky130_fd_pr__pfet_01v8 w=84 l=30
X23 Q a_1059_315# VGND VNB sky130_fd_pr__nfet_01v8 w=130 l=30
C0 a_27_47# a_466_413# 0.63fF
C1 a_27_47# D 0.21fF
C2 CLK D 0.05fF
C3 a_891_413# a_975_413# 0.05fF
C4 a_592_47# a_466_413# 0.02fF
C5 a_27_47# a_381_47# 0.21fF
C6 a_193_47# a_466_413# 0.38fF
C7 a_27_47# a_891_413# 0.09fF
C8 a_193_47# D 0.42fF
C9 CLK a_381_47# 0.02fF
C10 Q a_1059_315# 0.28fF
C11 a_466_413# VPB 0.01fF
C12 D VPB 0.00fF
C13 a_193_47# a_381_47# 0.26fF
C14 a_634_159# a_1059_315# 0.04fF
C15 a_193_47# a_891_413# 0.44fF
C16 VGND a_466_413# 0.17fF
C17 VGND D 0.06fF
C18 a_1059_315# VPWR 0.41fF
C19 a_381_47# VPB 0.00fF
C20 Q VPWR 0.23fF
C21 a_891_413# VPB 0.00fF
C22 VGND a_381_47# 0.11fF
C23 a_634_159# VPWR 0.23fF
C24 VGND a_891_413# 0.21fF
C25 D a_466_413# 0.04fF
C26 a_27_47# a_1059_315# 0.11fF
C27 a_561_413# VPWR 0.02fF
C28 a_466_413# a_381_47# 0.11fF
C29 D a_381_47# 0.35fF
C30 a_466_413# a_891_413# 0.03fF
C31 VPWR a_975_413# 0.02fF
C32 a_27_47# a_634_159# 0.37fF
C33 VGND a_1017_47# 0.01fF
C34 a_193_47# a_1059_315# 0.11fF
C35 a_27_47# VPWR 0.76fF
C36 a_193_47# Q 0.01fF
C37 CLK VPWR 0.06fF
C38 a_193_47# a_634_159# 0.28fF
C39 a_1059_315# VPB 0.01fF
C40 VGND a_1059_315# 0.26fF
C41 a_193_47# VPWR 0.42fF
C42 Q VPB 0.00fF
C43 a_634_159# VPB 0.00fF
C44 VGND Q 0.15fF
C45 a_634_159# VGND 0.26fF
C46 VPB VPWR 0.09fF
C47 VGND VPWR 0.03fF
C48 a_27_47# CLK 0.41fF
C49 a_1017_47# a_891_413# 0.04fF
C50 a_466_413# a_1059_315# 0.02fF
C51 a_193_47# a_27_47# 2.23fF
C52 a_193_47# CLK 0.06fF
C53 a_634_159# a_466_413# 0.59fF
C54 a_634_159# D 0.04fF
C55 a_27_47# VPB 0.01fF
C56 a_891_413# a_1059_315# 0.66fF
C57 a_466_413# VPWR 0.36fF
C58 D VPWR 0.03fF
C59 a_27_47# VGND 0.38fF
C60 Q a_891_413# 0.04fF
C61 CLK VPB 0.00fF
C62 a_634_159# a_381_47# 0.04fF
C63 a_466_413# a_561_413# 0.04fF
C64 a_634_159# a_891_413# 0.11fF
C65 VGND CLK 0.05fF
C66 a_193_47# VPB 0.01fF
C67 a_381_47# VPWR 0.14fF
C68 a_891_413# VPWR 0.22fF
C69 VGND a_592_47# 0.01fF
C70 a_193_47# VGND 0.29fF
C71 Q VNB 0.04fF
C72 VGND VNB 0.33fF
C73 VPWR VNB 0.35fF
C74 VPB VNB 0.29fF
C75 a_381_47# VNB 0.09fF
C76 a_891_413# VNB 0.39fF
C77 a_1059_315# VNB 0.58fF
C78 a_466_413# VNB 0.33fF
C79 a_634_159# VNB 0.35fF
C80 a_193_47# VNB 0.16fF
C81 a_27_47# VNB 0.34fF
.ends
