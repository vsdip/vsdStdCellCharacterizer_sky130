
    .include sky130nm.lib
    * /home/saurabh/esim-workspace/cmos_nand_gate/cmos_nand_gate.cir
* .include sky130nm.lib
.include example/esim/rahul_abskl.com_nitk/Half_Adder/xor.sub
.include example/esim/rahul_abskl.com_nitk/Half_Adder/and.sub
v1  A gnd pulse(0 1.8 0 0 0 17m 33m)
v2  B gnd pulse(0 1.8 0 0 0 10m 20m)
vc  vcc gnd dc 1.8
* u2  inputb plot_v1
* u1  inputa plot_v1
* u3  out plot_v1
x1 A B sum vcc xor
x2 A B cout vcc and
* .tran 0.1e-03 100e-03 0e-00

* Control Statements 

    CLOAD cout 0 1f
    .control
    let run  = 0 
 
    shell rm example/esim/rahul_abskl.com_nitk/Half_Adder/data/input_transition.txt
    shell rm example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_fall.txt
    shell rm example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_rise.txt
    shell rm example/esim/rahul_abskl.com_nitk/Half_Adder/data/fall_transition.txt
    shell rm example/esim/rahul_abskl.com_nitk/Half_Adder/data/rise_transition.txt
    foreach in_delay 0.01n 0.023n 0.0531329n 0.122474n 0.282311n 0.650743n 1.5n
    * Initiating Text Files in folder data
    echo "input_transition:$in_delay" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/input_transition.txt
    echo "input_transition:$in_delay" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_fall.txt
    echo "input_transition:$in_delay" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_rise.txt
    echo "input_transition:$in_delay" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/fall_transition.txt
    echo "input_transition:$in_delay" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/rise_transition.txt
    * 1.666 to match the slew rate
    let actual_rtime = $in_delay*1.666   

    * Input Vector - Load Cap values(index2)
    foreach out_cap 0.0005000000p 0.0012632050p 0.0031913740p 0.0080627180p 0.0203697300p 0.0514622900p 0.1300148000p
        reset
        
        * Changing the V2 Supply Rise time as per the Input Rise Time vector
        alter @v1[pulse] = [ 0 1.8 0 $&actual_rtime $&actual_rtime 50ns 100ns ]
        alter @v2[PWL] = [ 0 1.8 ]
        * Changing the C1 value as per the foreach list
        alter CLOAD $out_cap
        
        tran 0.01n 300ns
        run

        reset
        * Verification of INPUT RISE TIME
        meas tran ts1 when v(A)=1.4400000000000002 RISE=1 
        meas tran ts2 when v(A)=0.36000000000000004 RISE=1
        meas tran ts3 when v(A)=1.4400000000000002 FALL=1 
        meas tran ts4 when v(A)=0.36000000000000004 FALL=1
        let RISE_IN_SLEW = (ts1-ts2)/1n
        let FALL_IN_SLEW = (ts4-ts3)/1n
        echo "actual_rise_slew:$&RISE_IN_SLEW" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/input_transition.txt
        echo "actual_fall_slew:$&FALL_IN_SLEW" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/input_transition.txt


        print run
        * Measuring Cell Fall Time @ 50% of VDD(1.8V) 
        meas tran tinfall when v(A)=0.9 FALL=1 
        meas tran tofall when v(cout)=0.9 FALL=1
        let cfall = (tofall-tinfall)/1n
        if abs(cfall)>20
            meas tran tinfall when v(A)=0.9 Rise=1 
            meas tran tofall when v(cout)=0.9 FALL=1
            let cfall = abs(tofall-tinfall)/1n
        end
        print cfall
        echo "out_cap:$out_cap:cell_fall:$&cfall" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_fall.txt

        * Measuring Cell Rise Time @ 50% of VDD(1.8V) 
        meas tran tinrise when v(A)=0.9 RISE=1 
        meas tran torise when v(cout)=0.9 RISE=1
        let crise = (torise-tinrise)/1n
        if abs(crise)>20
            meas tran tinrise when v(A)=0.9 FALL=1 
            meas tran torise when v(cout)=0.9 RISE=1
            let crise = abs(tinrise-torise)/1n
        end
        print crise
        echo "out_cap:$out_cap:cell_rise:$&crise" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/cell_rise.txt

        * Measuring Fall transition Time @ 80-20% of VDD(1.8V) 
        meas tran ft1 when v(cout)=1.4400000000000002 FALL=2 
        meas tran ft2 when v(cout)=0.36000000000000004 FALL=2
        let fall_tran = (ft2-ft1)/1n
        print fall_tran
        echo "out_cap:$out_cap:fall_transition:$&fall_tran" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/fall_transition.txt
        
        * Measuring Rise transition Time @ 20-80% of VDD(1.8V) 
        meas tran rt1 when v(cout)=1.4400000000000002 RISE=2 
        meas tran rt2 when v(cout)=0.36000000000000004 RISE=2
        let rise_tran = ((rt1-rt2)/1n)
        print rise_tran
        echo "out_cap:$out_cap:rise_transition:$&rise_tran" >> example/esim/rahul_abskl.com_nitk/Half_Adder/data/rise_transition.txt
        let run = run + 1
        * plot a y
    end
    end
    quit
    .endc